localparam CLK_PERIOD           = 10;           // 10ns, 100MHz

localparam IMEM_WORD            = 4 * 1024;     // 16KB
localparam DMEM_WORD            = 16 * 1024;    // 64KB