timeunit 1ns;
timeprecision 1ps;

package uart_defines;
    `include "uart_parameter.svh"
    `include "uart_signal.svh"
endpackage